`timescale 1ns / 1ps

module mul_normalizer (
  input  [ 4:0] exponent,
  input  [21:0] mantissa_prod,
  output [14:0] result
);

  wire [4:0] result_exponent;
  wire [9:0] result_mantissa;

  assign result_exponent = (mantissa_prod[21]) ? (exponent + 1'b1): exponent;
  assign result_mantissa = (mantissa_prod[21]) ? mantissa_prod[20:11]:mantissa_prod[19:10];
  assign result          = {result_exponent,result_mantissa};

// No rounding and No overflow/underflow detection

endmodule
